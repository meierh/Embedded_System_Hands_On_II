package DCT;

interface DCT;
// Add custom interface definitions
endinterface

module mkDCT(DCT);

    rule doNothing;
        $display("Hello World!");
    endrule

endmodule

endpackage
